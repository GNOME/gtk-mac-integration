�� / *   W i n d o w s | B r i n g   A l l   T o   F r o n t   m e n u   i t e m   t i t l e   * / 
 " B r i n g   A l l   t o   F r o n t "   =   " T a   m e d   a l l a   l � n g s t   f r a m " ; 
 
 / *   H i d e   m e n u   i t e m   t i t l e   * / 
 " H i d e "   =   " D � l j " ; 
 
 / *   H i d e   O t h e r s   m e n u   i t e m   t i t l e   * / 
 " H i d e   O t h e r s "   =   " D � l j   m . f l . " ; 
 
 / *   W i n d o w s | M i n i m i z e   m e n u   i t e m   * / 
 " M i n i m i z e "   =   " M i n i m e r a " ; 
 
 / *   Q u i t   m e n u   i t e m   t i t l e   * / 
 " Q u i t "   =   " A v s l u t a " ; 
 
 / *   S e r v i c e s   M e n u   I t e m   t i t l e   * / 
 " S e r v i c e s "   =   " T j � n s t e r " ; 
 
 / *   S h o w   A l l   m e n u   i t e m   t i t l e   * / 
 " S h o w   A l l "   =   " V i s a   a l l a " ; 
 
 / *   W i n d o w   M e n u   t i t l e   * / 
 " W i n d o w "   =   " F � n s t e r " ; 
 
 / *   H e l p   M e n u   t i t l e   * / 
 " H e l p "   =   " H j � l p " ; 
